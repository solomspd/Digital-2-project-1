*** SPICE deck for cell NOR3_S1_simNEW{lay} from library NOR3
*** Created on Sun Apr 12, 2020 03:42:53
*** Last revised on Sun Apr 12, 2020 03:56:41
*** Written on Sun Apr 12, 2020 03:56:47 by Electric VLSI Design System, version 9.07
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF

*** SUBCIRCUIT NOR3__NOR3_S1 FROM CELL NOR3_S1{lay}
.SUBCKT NOR3__NOR3_S1 A B C gnd out vdd
Mnmos@0 gnd A out gnd NMOS L=0.36U W=0.9U AS=2.956P AD=2.997P PS=6.48U PD=8.46U
Mnmos@1 out B gnd gnd NMOS L=0.36U W=0.9U AS=2.997P AD=2.956P PS=8.46U PD=6.48U
Mnmos@2 gnd C out gnd NMOS L=0.36U W=0.9U AS=2.956P AD=2.997P PS=6.48U PD=8.46U
Mpmos@0 net@14 B net@13 vdd PMOS L=0.36U W=6.66U AS=3.742P AD=3.791P PS=14.4U PD=14.58U
Mpmos@3 net@13 C out vdd PMOS L=0.36U W=6.66U AS=2.956P AD=3.742P PS=6.48U PD=14.4U
Mpmos@4 vdd A net@14 vdd PMOS L=0.36U W=6.66U AS=3.791P AD=15.309P PS=14.58U PD=31.86U
.ENDS NOR3__NOR3_S1

*** TOP LEVEL CELL: NOR3_S1_simNEW{lay}
XNOR3_S1@0 IN_1 GND GND GND OUT VDD NOR3__NOR3_S1

* Spice Code nodes in cell cell 'NOR3_S1_simNEW{lay}'
vdd vdd 0 DC 3.3
vin IN_1 0 dc pulse 0 3.3 10n 667ps 667ps 10n
.tran 0 30n
cload OUT 0 53.16fF
.measure tpdr trig v(IN_1) val=1.67 fall=1 TARG v(OUT) val=1.67 rise=1
.measure tpdf trig v(IN_1) val=1.67 rise=1 TARG v(OUT) val=1.67 fall=1
.measure trise trig v(OUT) val=1 rise=1 TARG v(OUT) val=3.3 rise=1
.measure tfall trig v(OUT) val=3.3 fall=1 TARG v(OUT) val=1 fall=1
.include C:\Electric\scmos18.txt
.END
.END
