*** SPICE deck for cell somp_sim_lay{lay} from library test1
*** Created on Sun Apr 05, 2020 06:26:11
*** Last revised on Tue Apr 14, 2020 05:33:33
*** Written on Tue Apr 14, 2020 05:34:11 by Electric VLSI Design System, version 9.07
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF

*** SUBCIRCUIT test1__comp FROM CELL comp{lay}
.SUBCKT test1__comp F gnd vdd W X Z
Mnmos@0 net@29 X gnd gnd NMOS L=0.36U W=0.9U AS=3.888P AD=0.486P PS=11.34U PD=1.98U
Mnmos@1 F net@39 net@29 gnd N L=0.36U W=0.9U AS=0.486P AD=1.223P PS=1.98U PD=3.96U
Mnmos@2 net@30 W F gnd N L=0.36U W=0.9U AS=1.223P AD=0.486P PS=3.96U PD=1.98U
Mnmos@3 gnd Z net@30 gnd N L=0.36U W=0.9U AS=0.486P AD=3.888P PS=1.98U PD=11.34U
Mpmos@1 net@4 net@39 vdd vdd P L=0.36U W=1.98U AS=4.714P AD=1.366P PS=12.06U PD=4.02U
Mpmos@2 net@4 W F vdd P L=0.36U W=1.98U AS=1.223P AD=1.366P PS=3.96U PD=4.02U
Mpmos@3 F Z net@4 vdd PMOS L=0.36U W=1.98U AS=1.366P AD=1.223P PS=4.02U PD=3.96U
Mpmos@4 vdd X net@36 vdd P L=0.36U W=1.98U AS=1.96P AD=4.714P PS=5.94U PD=12.06U
.ENDS test1__comp

*** TOP LEVEL CELL: somp_sim_lay{lay}
Xcomp@0 F comp@0_GND comp@0_VDD W X Z test1__comp

* Spice Code nodes in cell cell 'somp_sim_lay{lay}'
.param transsi=166.66p
vdd VDD 0 DC 3.3
vw W 0 pulse 3.3 0 1u {transsi} {transsi} 2u 4u
vx X 0 DC 3.3
vy Y 0 DC 3.3
vz Z 0 DC 3.3
*vx X 0 pulse 3.3 0 0 {transsi} {transsi} 0u 10u
*vy Y 0 pulse 3.3 0 0 {transsi} {transsi} 0u 10u
*vz Z 0 pulse 3.3 0 0 {transsi} {transsi} 0u 10u
cload F 0 26.58fF
.tran 0 10u
.measure tdpr trig v(W) val=1.65 fall =1 TARG v(F) val=1.65 rise=1
.measure tdpf trig v(W) val=1.65 rise =1 TARG v(F) val=1.65 fall=1
.measure trise trig v(F) val=0.66 rise =1 TARG v(F) val=2.64 rise=1
.measure tfall trig v(F) val=2.64 fall =1 TARG v(F) val=0.66 fall=1
.include '/data/Abdo/Abdo/Abdo's University work/spring 2020/Digital 2/Project1/Digital-2-project-1/scmos18(2).txt'
.END
