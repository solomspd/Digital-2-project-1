*** SPICE deck for cell comp_sz8_sim{lay} from library test1
*** Created on Tue Apr 14, 2020 06:56:28
*** Last revised on Tue Apr 14, 2020 07:02:14
*** Written on Tue Apr 14, 2020 07:03:18 by Electric VLSI Design System, version 9.07
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF

*** SUBCIRCUIT test1__comp_sz8 FROM CELL comp_sz8{lay}
.SUBCKT test1__comp_sz8 F gnd vdd W X Y Z
Mnmos@0 net@1 X gnd gnd NMOS L=0.36U W=7.2U AS=10.125P AD=3.888P PS=23.94U PD=8.28U
Mnmos@1 F Y net@1 gnd N L=0.36U W=7.2U AS=3.888P AD=9.785P PS=8.28U PD=20.97U
Mnmos@2 net@13 W F gnd N L=0.36U W=7.2U AS=9.785P AD=3.888P PS=20.97U PD=8.28U
Mnmos@3 gnd Z net@13 gnd N L=0.36U W=7.2U AS=3.888P AD=10.125P PS=8.28U PD=23.94U
Mpmos@0 vdd X net@5 vdd PMOS L=0.36U W=15.84U AS=12.118P AD=12.199P PS=25.29U PD=25.92U
Mpmos@1 net@5 Y vdd vdd P L=0.36U W=15.84U AS=12.199P AD=12.118P PS=25.92U PD=25.29U
Mpmos@2 net@5 W F vdd P L=0.36U W=15.84U AS=9.785P AD=12.118P PS=20.97U PD=25.29U
Mpmos@3 F Z net@5 vdd P L=0.36U W=15.84U AS=12.118P AD=9.785P PS=25.29U PD=20.97U
.ENDS test1__comp_sz8

*** TOP LEVEL CELL: comp_sz8_sim{lay}
Xcomp_sz8@0 F GND VDD W X Y Z test1__comp_sz8

* Spice Code nodes in cell cell 'comp_sz8_sim{lay}'
.param transsi=1333.33p
vdd VDD 0 DC 3.3
vw W 0 pulse 3.3 0 1u {transsi} {transsi} 2u 4u
vx X 0 DC 3.3
vy Y 0 DC 0
vz Z 0 DC 3.3
*vx X 0 pulse 3.3 0 0 {transsi} {transsi} 0u 10u
*vy Y 0 pulse 3.3 0 0 {transsi} {transsi} 0u 10u
*vz Z 0 pulse 3.3 0 0 {transsi} {transsi} 0u 10u
cload F 0 1333.33fF
.tran 0 10u
.measure tdpr trig v(W) val=1.65 fall =1 TARG v(F) val=1.65 rise=1
.measure tdpf trig v(W) val=1.65 rise =1 TARG v(F) val=1.65 fall=1
.measure trise trig v(F) val=0.66 rise =1 TARG v(F) val=2.64 rise=1
.measure tfall trig v(F) val=2.64 fall =1 TARG v(F) val=0.66 fall=1
.include '/data/Abdo/Abdo/Abdo's University work/spring 2020/Digital 2/Project1/Digital-2-project-1/scmos18(2).txt'
.END
