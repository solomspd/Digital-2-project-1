*** SPICE deck for cell comp_sz2_sim{lay} from library test1
*** Created on Mon Apr 13, 2020 22:14:22
*** Last revised on Tue Apr 14, 2020 07:02:30
*** Written on Tue Apr 14, 2020 07:21:13 by Electric VLSI Design System, version 9.07
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF

*** SUBCIRCUIT test1__comp_sz2 FROM CELL comp_sz2{lay}
.SUBCKT test1__comp_sz2 F gnd vdd W X Y Z
Mnmos@4 net@1 X gnd gnd NMOS L=0.36U W=1.8U AS=4.779P AD=0.972P PS=13.14U PD=2.88U
Mnmos@5 F Y net@1 gnd N L=0.36U W=1.8U AS=0.972P AD=2.446P PS=2.88U PD=6.39U
Mnmos@6 net@4 W F gnd N L=0.36U W=1.8U AS=2.446P AD=0.972P PS=6.39U PD=2.88U
Mnmos@7 gnd Z net@4 gnd N L=0.36U W=1.8U AS=0.972P AD=4.779P PS=2.88U PD=13.14U
Mpmos@0 vdd X net@6 vdd PMOS L=0.36U W=3.96U AS=3.029P AD=5.783P PS=7.47U PD=14.04U
Mpmos@1 net@6 Y vdd vdd P L=0.36U W=3.96U AS=5.783P AD=3.029P PS=14.04U PD=7.47U
Mpmos@2 net@6 W F vdd P L=0.36U W=3.96U AS=2.446P AD=3.029P PS=6.39U PD=7.47U
Mpmos@3 F Z net@6 vdd P L=0.36U W=3.96U AS=3.029P AD=2.446P PS=7.47U PD=6.39U
.ENDS test1__comp_sz2

*** TOP LEVEL CELL: comp_sz2_sim{lay}
Xcomp_sz2@1 F GND VDD W X Y Z test1__comp_sz2

* Spice Code nodes in cell cell 'comp_sz2_sim{lay}'
.param transsi=166.66p
vdd VDD 0 DC 3.3
vw W 0 pulse 3.3 0 1u {transsi} {transsi} 2u 4u
vx X 0 DC 3.3
vy Y 0 DC 0
vz Z 0 DC 3.3
*vx X 0 pulse 3.3 0 0 {transsi} {transsi} 0u 10u
*vy Y 0 pulse 3.3 0 0 {transsi} {transsi} 0u 10u
*vz Z 0 pulse 3.3 0 0 {transsi} {transsi} 0u 10u
cload F 0 26.58fF
.tran 0 10u
.measure tdpr trig v(W) val=1.65 fall =1 TARG v(F) val=1.65 rise=1
.measure tdpf trig v(W) val=1.65 rise =1 TARG v(F) val=1.65 fall=1
.measure trise trig v(F) val=0.66 rise =1 TARG v(F) val=2.64 rise=1
.measure tfall trig v(F) val=2.64 fall =1 TARG v(F) val=0.66 fall=1
.include '/data/Abdo/Abdo/Abdo's University work/spring 2020/Digital 2/Project1/Digital-2-project-1/scmos18(2).txt'
.END
