*** SPICE deck for cell somp_sim_lay{lay} from library noname
*** Created on Sun Apr 05, 2020 06:26:11
*** Last revised on Sun Apr 12, 2020 18:05:03
*** Written on Sun Apr 12, 2020 18:06:09 by Electric VLSI Design System, version 9.07
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF

*** SUBCIRCUIT noname__comp FROM CELL noname:comp{lay}
.SUBCKT noname__comp gnd out vdd W X Y Z
Mnmos@0 net@29 Y gnd gnd NMOS L=0.36U W=0.9U AS=4.739P AD=0.535P PS=13.23U PD=2.52U
Mnmos@1 out Z net@29 gnd N L=0.36U W=0.9U AS=0.535P AD=1.867P PS=2.52U PD=5.445U
Mnmos@2 net@30 W out gnd N L=0.36U W=0.9U AS=1.867P AD=0.583P PS=5.445U PD=2.7U
Mnmos@3 gnd X net@30 gnd N L=0.36U W=0.9U AS=0.583P AD=4.739P PS=2.7U PD=13.23U
Mpmos@0 vdd Y net@2 vdd P L=0.36U W=2.16U AS=1.993P AD=5.411P PS=5.085U PD=13.32U
Mpmos@1 net@2 Z vdd vdd P L=0.36U W=2.16U AS=5.411P AD=1.993P PS=13.32U PD=5.085U
Mpmos@2 net@2 W out vdd P L=0.36U W=2.16U AS=1.867P AD=1.993P PS=5.445U PD=5.085U
Mpmos@3 out X net@2 vdd PMOS L=0.36U W=2.16U AS=1.993P AD=1.867P PS=5.085U PD=5.445U
.ENDS noname__comp

*** TOP LEVEL CELL: noname:somp_sim_lay{lay}
Xcomp@0 GND F VDD W X Y Z noname__comp

.param transsi=166.66p

* Spice Code nodes in cell cell 'noname:somp_sim_lay{lay}'
vdd VDD 0 DC 3.3
vw W 0 pulse 3.3 0 0 {transsi} {transsi} 1u 2u
vx X 0 pulse 3.3 0 0 {transsi} {transsi} 2u 4u
vy Y 0 pulse 3.3 0 0 {transsi} {transsi} 4u 8u
vz Z 0 pulse 3.3 0 0 {transsi} {transsi} 8u 16u
cload F 0 13.29fF
.tran 0 10u
.measure tdpr trig v(W) val=1.65 fall =1 TARG v(F) val=1.65 rise=1
.measure tdpf trig v(W) val=1.65 rise =1 TARG v(F) val=1.65 fall=1
.measure trise trig v(F) val=0.66 rise =1 TARG v(F) val=2.64 rise=1
.measure tfall trig v(F) val=2.64 fall =1 TARG v(F) val=0.66 fall=1
.include '/data/Abdo/Abdo/Abdo's University work/spring 2020/Digital 2/Project1/Digital-2-project-1/scmos18(2).txt'
.END
